-------------------------------------
-- Defines the dataPath width
--
-------------------------------------
package mypackage is
   constant XBITS :INTEGER := 8; 
   constant YBITS :INTEGER := 8;
   constant GRAIN :INTEGER := 2; --Allways in 2!!!!
end mypackage;
